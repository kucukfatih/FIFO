`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.03.2024 22:54:57
// Design Name: 
// Module Name: comp
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module comp#(parameter K = 3)(

input wire [K-1:0] A,B,
output wire equal_flag,
output wire zero_flag

    );
    
assign equal_flag = (A == B) ? 1'b1 : 1'b0;

assign zero_flag = (B == 0) ? 1'b1 : 1'b0;

endmodule
